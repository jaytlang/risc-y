// `define MEM_LAT 10
