import RegFile::*;
import BRAM::*;
