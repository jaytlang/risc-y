// Copyright (c) 2017 Massachusetts Institute of Technology
//
// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

import BRAMCore::*;
import FIFOF::*;
import SpecialFIFOs::*;

interface RWBramCore#(type addrT, type dataT);
   method Action wrReq(addrT a, dataT d);
   method Action rdReq(addrT a);
   method dataT rdResp;
   method Bool rdRespValid;
   method Action deqRdResp;
endinterface

module mkRWBramCore(RWBramCore#(addrT, dataT)) provisos(
   Bits#(addrT, addrSz), Bits#(dataT, dataSz)
   );
   BRAM_DUAL_PORT#(addrT, dataT) bram <- mkBRAMCore2(valueOf(TExp#(addrSz)), False);
   BRAM_PORT#(addrT, dataT) wrPort = bram.a;
   BRAM_PORT#(addrT, dataT) rdPort = bram.b;
   
   // 1 elem pipeline fifo to add guard for read req/resp
   // must be 1 elem to make sure rdResp is not corrupted
   // BRAMCore should not change output if no req is made
   FIFOF#(void) rdReqQ <- mkPipelineFIFOF;
   
   method Action wrReq(addrT a, dataT d);
      wrPort.put(True, a, d);
   endmethod
   
   method Action rdReq(addrT a);
      rdReqQ.enq(?);
      rdPort.put(False, a, ?);
   endmethod
   
   method dataT rdResp if(rdReqQ.notEmpty);
      return rdPort.read;
   endmethod
   
   method rdRespValid = rdReqQ.notEmpty;
   
   method Action deqRdResp;
      rdReqQ.deq;
   endmethod
endmodule
